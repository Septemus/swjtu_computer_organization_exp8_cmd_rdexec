library verilog;
use verilog.vl_types.all;
entity exp8_vlg_vec_tst is
end exp8_vlg_vec_tst;
